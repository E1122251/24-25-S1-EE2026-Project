`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 10/20/2024 06:09:59 PM
// Design Name: 
// Module Name: screen_after_collision
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module screen_after_collision(
    input clock_100mhz,
    input [12:0] pixel_index,
    input game_active,
    input is_collision,
    input btnC,
    
    output reg [15:0] oled_data_collision,
    output reg return_to_menu = 0
    );
    reg [31:0] count = 0;
    always @ (posedge clock_100mhz)begin
        if (game_active==0) begin
            return_to_menu <= 0;
            count <= 0;
        end
        if (game_active==1 && is_collision==1) begin
            if (count == 32'd100_000_000) begin
                if (btnC == 1) begin
                    return_to_menu <= 1 ; // 
                    count <= 0;
                    end
                else begin
                    count <= count;
                    end
                end
            else begin
                count <= count +1;
                end
        end
    end
    
    
    //xy coordinate
    wire [6:0] x = pixel_index % 96;
    wire [5:0] y = pixel_index / 96;
    
    //for circle
    wire signed [8:0] dx = $signed({1'b0,x})-54;  //x-center 48
    wire signed [8:0] dy = $signed({1'b0,y})-73; //handle top from base 25, circle size 61, thickness 5 
    wire [16:0] square_dx = dx*dx;
    wire [16:0] square_dy = dy*dy;    
    wire [16:0] square_distance = square_dx + square_dy;
    
    always @ (posedge clock_100mhz)begin
        if (square_distance >= 900 && square_distance <= 1225) begin //handle
             oled_data_collision <= 16'hFD20; //orange
             end
        else if ((x >= 24 && x <= 96) && (y >=45  && y <= 48)) begin //grey line of insde car
                 oled_data_collision <= 16'h4929; // grey
                 end
        else if (y >= (51 - (x-18)) && //triangle at the end of grey line
                y <= (51 - (10 * (x-18) / 20)) &&  
                x >= 18 && x <= 24 // 
                )begin
                oled_data_collision <= 16'h4929;
                end 
        else if ((x >= 18 && x <= 96) && (y >= 42 && y <= 64)) begin //black square bottom (car display)
            oled_data_collision <= 16'h0000;
            end
            //17 44
            //11 43
        //using trapesium calculation to draw window frame
        else if (x <= (22 + (10 * y) / 40) && // right slent of trapezium 
            x >= (4 + (10 * y) / 30) &&  //left slent of trapezium, every increasement of y will cause x to be increase by 1/3
            y >= 0 && y <= 43 // 
            )begin
            oled_data_collision <= 16'h0000;
            end
        else if (x <= (96 - (11 * (y-6))) && //top window frame
            x >= (0 + (10 * (y-6)) / 10) &&  
            y >= 6 && y <= 13 // 
            )begin
            oled_data_collision <= 16'h0000;
            end
        else if ((x >= 0 && x <= 96) && (y >= 0 && y <= 6)) begin//top window frame square
                oled_data_collision <= 16'h000;
            end
        else if (y >= (53 - (10 * x) / 20) && //left window frame
            y <= 64 &&  
            x >= 0 && x <= 19 // 
            )begin
            oled_data_collision <= 16'h0000;
            end
        else if ((x >= 0 && x <= 8) && (y >= 46 && y <= 51)) begin//side miirror mirror
            oled_data_collision <= 16'h001F;
            end
        else if (x <= (9 + (10 * (y-42)) / 10) && //side mirror frame
            x >= 0 &&  
            y >= 42 && y <= 64 // 
            )begin
            oled_data_collision <= 16'h4929;
            end      
        else begin
            oled_data_collision <= 16'h83DD; //skyblue
        end
    end
    
    
    
endmodule
